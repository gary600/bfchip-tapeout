// THIS FILE IS OVERWRITTEN BY THE BUILD PIPELINE
module dummy;
	generate
		$error("chip.sv was not overwritten by the build pipeline");
	endgenerate
endmodule